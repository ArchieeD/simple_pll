magic
tech sky130A
magscale 1 2
timestamp 1741065640
<< nwell >>
rect -101 261 2804 582
<< pwell >>
rect 29 -17 63 17
rect 444 -17 478 17
rect 859 -17 893 17
rect 1274 -17 1308 17
rect 1689 -17 1723 17
rect 2104 -17 2138 17
rect 2519 -17 2553 17
<< scnmos >>
rect 120 47 150 177
rect 535 47 565 177
rect 950 47 980 177
rect 1365 47 1395 177
rect 1780 47 1810 177
rect 2195 47 2225 177
rect 2610 47 2640 177
<< scpmoshvt >>
rect 120 297 150 497
rect 535 297 565 497
rect 950 297 980 497
rect 1365 297 1395 497
rect 1780 297 1810 497
rect 2195 297 2225 497
rect 2610 297 2640 497
<< ndiff >>
rect 68 165 120 177
rect 68 131 76 165
rect 110 131 120 165
rect 68 97 120 131
rect 68 63 76 97
rect 110 63 120 97
rect 68 47 120 63
rect 150 165 202 177
rect 150 131 160 165
rect 194 131 202 165
rect 150 97 202 131
rect 150 63 160 97
rect 194 63 202 97
rect 150 47 202 63
rect 483 165 535 177
rect 483 131 491 165
rect 525 131 535 165
rect 483 97 535 131
rect 483 63 491 97
rect 525 63 535 97
rect 483 47 535 63
rect 565 165 617 177
rect 565 131 575 165
rect 609 131 617 165
rect 565 97 617 131
rect 565 63 575 97
rect 609 63 617 97
rect 565 47 617 63
rect 898 165 950 177
rect 898 131 906 165
rect 940 131 950 165
rect 898 97 950 131
rect 898 63 906 97
rect 940 63 950 97
rect 898 47 950 63
rect 980 165 1032 177
rect 980 131 990 165
rect 1024 131 1032 165
rect 980 97 1032 131
rect 980 63 990 97
rect 1024 63 1032 97
rect 980 47 1032 63
rect 1313 165 1365 177
rect 1313 131 1321 165
rect 1355 131 1365 165
rect 1313 97 1365 131
rect 1313 63 1321 97
rect 1355 63 1365 97
rect 1313 47 1365 63
rect 1395 165 1447 177
rect 1395 131 1405 165
rect 1439 131 1447 165
rect 1395 97 1447 131
rect 1395 63 1405 97
rect 1439 63 1447 97
rect 1395 47 1447 63
rect 1728 165 1780 177
rect 1728 131 1736 165
rect 1770 131 1780 165
rect 1728 97 1780 131
rect 1728 63 1736 97
rect 1770 63 1780 97
rect 1728 47 1780 63
rect 1810 165 1862 177
rect 1810 131 1820 165
rect 1854 131 1862 165
rect 1810 97 1862 131
rect 1810 63 1820 97
rect 1854 63 1862 97
rect 1810 47 1862 63
rect 2143 165 2195 177
rect 2143 131 2151 165
rect 2185 131 2195 165
rect 2143 97 2195 131
rect 2143 63 2151 97
rect 2185 63 2195 97
rect 2143 47 2195 63
rect 2225 165 2277 177
rect 2225 131 2235 165
rect 2269 131 2277 165
rect 2225 97 2277 131
rect 2225 63 2235 97
rect 2269 63 2277 97
rect 2225 47 2277 63
rect 2558 165 2610 177
rect 2558 131 2566 165
rect 2600 131 2610 165
rect 2558 97 2610 131
rect 2558 63 2566 97
rect 2600 63 2610 97
rect 2558 47 2610 63
rect 2640 165 2692 177
rect 2640 131 2650 165
rect 2684 131 2692 165
rect 2640 97 2692 131
rect 2640 63 2650 97
rect 2684 63 2692 97
rect 2640 47 2692 63
<< pdiff >>
rect 68 485 120 497
rect 68 451 76 485
rect 110 451 120 485
rect 68 417 120 451
rect 68 383 76 417
rect 110 383 120 417
rect 68 349 120 383
rect 68 315 76 349
rect 110 315 120 349
rect 68 297 120 315
rect 150 485 202 497
rect 150 451 160 485
rect 194 451 202 485
rect 483 485 535 497
rect 150 417 202 451
rect 150 383 160 417
rect 194 383 202 417
rect 150 349 202 383
rect 150 315 160 349
rect 194 315 202 349
rect 483 451 491 485
rect 525 451 535 485
rect 483 417 535 451
rect 483 383 491 417
rect 525 383 535 417
rect 483 349 535 383
rect 150 297 202 315
rect 483 315 491 349
rect 525 315 535 349
rect 483 297 535 315
rect 565 485 617 497
rect 565 451 575 485
rect 609 451 617 485
rect 898 485 950 497
rect 565 417 617 451
rect 565 383 575 417
rect 609 383 617 417
rect 565 349 617 383
rect 565 315 575 349
rect 609 315 617 349
rect 898 451 906 485
rect 940 451 950 485
rect 898 417 950 451
rect 898 383 906 417
rect 940 383 950 417
rect 898 349 950 383
rect 565 297 617 315
rect 898 315 906 349
rect 940 315 950 349
rect 898 297 950 315
rect 980 485 1032 497
rect 980 451 990 485
rect 1024 451 1032 485
rect 1313 485 1365 497
rect 980 417 1032 451
rect 980 383 990 417
rect 1024 383 1032 417
rect 980 349 1032 383
rect 980 315 990 349
rect 1024 315 1032 349
rect 1313 451 1321 485
rect 1355 451 1365 485
rect 1313 417 1365 451
rect 1313 383 1321 417
rect 1355 383 1365 417
rect 1313 349 1365 383
rect 980 297 1032 315
rect 1313 315 1321 349
rect 1355 315 1365 349
rect 1313 297 1365 315
rect 1395 485 1447 497
rect 1395 451 1405 485
rect 1439 451 1447 485
rect 1728 485 1780 497
rect 1395 417 1447 451
rect 1395 383 1405 417
rect 1439 383 1447 417
rect 1395 349 1447 383
rect 1395 315 1405 349
rect 1439 315 1447 349
rect 1728 451 1736 485
rect 1770 451 1780 485
rect 1728 417 1780 451
rect 1728 383 1736 417
rect 1770 383 1780 417
rect 1728 349 1780 383
rect 1395 297 1447 315
rect 1728 315 1736 349
rect 1770 315 1780 349
rect 1728 297 1780 315
rect 1810 485 1862 497
rect 1810 451 1820 485
rect 1854 451 1862 485
rect 2143 485 2195 497
rect 1810 417 1862 451
rect 1810 383 1820 417
rect 1854 383 1862 417
rect 1810 349 1862 383
rect 1810 315 1820 349
rect 1854 315 1862 349
rect 2143 451 2151 485
rect 2185 451 2195 485
rect 2143 417 2195 451
rect 2143 383 2151 417
rect 2185 383 2195 417
rect 2143 349 2195 383
rect 1810 297 1862 315
rect 2143 315 2151 349
rect 2185 315 2195 349
rect 2143 297 2195 315
rect 2225 485 2277 497
rect 2225 451 2235 485
rect 2269 451 2277 485
rect 2558 485 2610 497
rect 2225 417 2277 451
rect 2225 383 2235 417
rect 2269 383 2277 417
rect 2225 349 2277 383
rect 2225 315 2235 349
rect 2269 315 2277 349
rect 2558 451 2566 485
rect 2600 451 2610 485
rect 2558 417 2610 451
rect 2558 383 2566 417
rect 2600 383 2610 417
rect 2558 349 2610 383
rect 2225 297 2277 315
rect 2558 315 2566 349
rect 2600 315 2610 349
rect 2558 297 2610 315
rect 2640 485 2692 497
rect 2640 451 2650 485
rect 2684 451 2692 485
rect 2640 417 2692 451
rect 2640 383 2650 417
rect 2684 383 2692 417
rect 2640 349 2692 383
rect 2640 315 2650 349
rect 2684 315 2692 349
rect 2640 297 2692 315
<< ndiffc >>
rect 76 131 110 165
rect 76 63 110 97
rect 160 131 194 165
rect 160 63 194 97
rect 491 131 525 165
rect 491 63 525 97
rect 575 131 609 165
rect 575 63 609 97
rect 906 131 940 165
rect 906 63 940 97
rect 990 131 1024 165
rect 990 63 1024 97
rect 1321 131 1355 165
rect 1321 63 1355 97
rect 1405 131 1439 165
rect 1405 63 1439 97
rect 1736 131 1770 165
rect 1736 63 1770 97
rect 1820 131 1854 165
rect 1820 63 1854 97
rect 2151 131 2185 165
rect 2151 63 2185 97
rect 2235 131 2269 165
rect 2235 63 2269 97
rect 2566 131 2600 165
rect 2566 63 2600 97
rect 2650 131 2684 165
rect 2650 63 2684 97
<< pdiffc >>
rect 76 451 110 485
rect 76 383 110 417
rect 76 315 110 349
rect 160 451 194 485
rect 160 383 194 417
rect 160 315 194 349
rect 491 451 525 485
rect 491 383 525 417
rect 491 315 525 349
rect 575 451 609 485
rect 575 383 609 417
rect 575 315 609 349
rect 906 451 940 485
rect 906 383 940 417
rect 906 315 940 349
rect 990 451 1024 485
rect 990 383 1024 417
rect 990 315 1024 349
rect 1321 451 1355 485
rect 1321 383 1355 417
rect 1321 315 1355 349
rect 1405 451 1439 485
rect 1405 383 1439 417
rect 1405 315 1439 349
rect 1736 451 1770 485
rect 1736 383 1770 417
rect 1736 315 1770 349
rect 1820 451 1854 485
rect 1820 383 1854 417
rect 1820 315 1854 349
rect 2151 451 2185 485
rect 2151 383 2185 417
rect 2151 315 2185 349
rect 2235 451 2269 485
rect 2235 383 2269 417
rect 2235 315 2269 349
rect 2566 451 2600 485
rect 2566 383 2600 417
rect 2566 315 2600 349
rect 2650 451 2684 485
rect 2650 383 2684 417
rect 2650 315 2684 349
<< psubdiff >>
rect -64 160 14 190
rect -64 81 -51 160
rect 1 81 14 160
rect -64 55 14 81
rect 351 160 429 190
rect 351 81 364 160
rect 416 81 429 160
rect 351 55 429 81
rect 766 160 844 190
rect 766 81 779 160
rect 831 81 844 160
rect 766 55 844 81
rect 1181 160 1259 190
rect 1181 81 1194 160
rect 1246 81 1259 160
rect 1181 55 1259 81
rect 1596 160 1674 190
rect 1596 81 1609 160
rect 1661 81 1674 160
rect 1596 55 1674 81
rect 2011 160 2089 190
rect 2011 81 2024 160
rect 2076 81 2089 160
rect 2011 55 2089 81
rect 2426 160 2504 190
rect 2426 81 2439 160
rect 2491 81 2504 160
rect 2426 55 2504 81
<< nsubdiff >>
rect -64 448 14 479
rect -64 385 -51 448
rect 3 385 14 448
rect -64 336 14 385
rect 351 448 429 479
rect 351 385 364 448
rect 418 385 429 448
rect 351 336 429 385
rect 766 448 844 479
rect 766 385 779 448
rect 833 385 844 448
rect 766 336 844 385
rect 1181 448 1259 479
rect 1181 385 1194 448
rect 1248 385 1259 448
rect 1181 336 1259 385
rect 1596 448 1674 479
rect 1596 385 1609 448
rect 1663 385 1674 448
rect 1596 336 1674 385
rect 2011 448 2089 479
rect 2011 385 2024 448
rect 2078 385 2089 448
rect 2011 336 2089 385
rect 2426 448 2504 479
rect 2426 385 2439 448
rect 2493 385 2504 448
rect 2426 336 2504 385
<< psubdiffcont >>
rect -51 81 1 160
rect 364 81 416 160
rect 779 81 831 160
rect 1194 81 1246 160
rect 1609 81 1661 160
rect 2024 81 2076 160
rect 2439 81 2491 160
<< nsubdiffcont >>
rect -51 385 3 448
rect 364 385 418 448
rect 779 385 833 448
rect 1194 385 1248 448
rect 1609 385 1663 448
rect 2024 385 2078 448
rect 2439 385 2493 448
<< poly >>
rect 120 497 150 523
rect 535 497 565 523
rect 950 497 980 523
rect 1365 497 1395 523
rect 1780 497 1810 523
rect 2195 497 2225 523
rect 2610 497 2640 523
rect 120 265 150 297
rect 535 265 565 297
rect 950 265 980 297
rect 1365 265 1395 297
rect 1780 265 1810 297
rect 2195 265 2225 297
rect 2610 265 2640 297
rect 64 249 150 265
rect 64 215 80 249
rect 114 215 150 249
rect 64 199 150 215
rect 479 249 565 265
rect 479 215 495 249
rect 529 215 565 249
rect 479 199 565 215
rect 894 249 980 265
rect 894 215 910 249
rect 944 215 980 249
rect 894 199 980 215
rect 1309 249 1395 265
rect 1309 215 1325 249
rect 1359 215 1395 249
rect 1309 199 1395 215
rect 1724 249 1810 265
rect 1724 215 1740 249
rect 1774 215 1810 249
rect 1724 199 1810 215
rect 2139 249 2225 265
rect 2139 215 2155 249
rect 2189 215 2225 249
rect 2139 199 2225 215
rect 2554 249 2640 265
rect 2554 215 2570 249
rect 2604 215 2640 249
rect 2554 199 2640 215
rect 120 177 150 199
rect 535 177 565 199
rect 950 177 980 199
rect 1365 177 1395 199
rect 1780 177 1810 199
rect 2195 177 2225 199
rect 2610 177 2640 199
rect 120 21 150 47
rect 535 21 565 47
rect 950 21 980 47
rect 1365 21 1395 47
rect 1780 21 1810 47
rect 2195 21 2225 47
rect 2610 21 2640 47
<< polycont >>
rect 80 215 114 249
rect 495 215 529 249
rect 910 215 944 249
rect 1325 215 1359 249
rect 1740 215 1774 249
rect 2155 215 2189 249
rect 2570 215 2604 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 415 527 444 561
rect 478 527 536 561
rect 570 527 628 561
rect 662 527 691 561
rect 830 527 859 561
rect 893 527 951 561
rect 985 527 1043 561
rect 1077 527 1106 561
rect 1245 527 1274 561
rect 1308 527 1366 561
rect 1400 527 1458 561
rect 1492 527 1521 561
rect 1660 527 1689 561
rect 1723 527 1781 561
rect 1815 527 1873 561
rect 1907 527 1936 561
rect 2075 527 2104 561
rect 2138 527 2196 561
rect 2230 527 2288 561
rect 2322 527 2351 561
rect 2490 527 2519 561
rect 2553 527 2611 561
rect 2645 527 2703 561
rect 2737 527 2766 561
rect 68 485 110 527
rect 68 466 76 485
rect -64 451 76 466
rect -64 448 110 451
rect -64 385 -51 448
rect 3 417 110 448
rect 3 385 76 417
rect -64 383 76 385
rect -64 359 110 383
rect 68 349 110 359
rect 68 315 76 349
rect 68 299 110 315
rect 144 485 210 493
rect 144 451 160 485
rect 194 451 210 485
rect 483 485 525 527
rect 483 466 491 485
rect 144 417 210 451
rect 144 383 160 417
rect 194 383 210 417
rect 144 349 210 383
rect 351 451 491 466
rect 351 448 525 451
rect 351 385 364 448
rect 418 417 525 448
rect 418 385 491 417
rect 351 383 491 385
rect 351 359 525 383
rect 144 315 160 349
rect 194 315 210 349
rect 144 297 210 315
rect 483 349 525 359
rect 483 315 491 349
rect 483 299 525 315
rect 559 485 625 493
rect 559 451 575 485
rect 609 451 625 485
rect 898 485 940 527
rect 898 466 906 485
rect 559 417 625 451
rect 559 383 575 417
rect 609 383 625 417
rect 559 349 625 383
rect 766 451 906 466
rect 766 448 940 451
rect 766 385 779 448
rect 833 417 940 448
rect 833 385 906 417
rect 766 383 906 385
rect 766 359 940 383
rect 559 315 575 349
rect 609 315 625 349
rect 559 297 625 315
rect 898 349 940 359
rect 898 315 906 349
rect 898 299 940 315
rect 974 485 1040 493
rect 974 451 990 485
rect 1024 451 1040 485
rect 1313 485 1355 527
rect 1313 466 1321 485
rect 974 417 1040 451
rect 974 383 990 417
rect 1024 383 1040 417
rect 974 349 1040 383
rect 1181 451 1321 466
rect 1181 448 1355 451
rect 1181 385 1194 448
rect 1248 417 1355 448
rect 1248 385 1321 417
rect 1181 383 1321 385
rect 1181 359 1355 383
rect 974 315 990 349
rect 1024 315 1040 349
rect 974 297 1040 315
rect 1313 349 1355 359
rect 1313 315 1321 349
rect 1313 299 1355 315
rect 1389 485 1455 493
rect 1389 451 1405 485
rect 1439 451 1455 485
rect 1728 485 1770 527
rect 1728 466 1736 485
rect 1389 417 1455 451
rect 1389 383 1405 417
rect 1439 383 1455 417
rect 1389 349 1455 383
rect 1596 451 1736 466
rect 1596 448 1770 451
rect 1596 385 1609 448
rect 1663 417 1770 448
rect 1663 385 1736 417
rect 1596 383 1736 385
rect 1596 359 1770 383
rect 1389 315 1405 349
rect 1439 315 1455 349
rect 1389 297 1455 315
rect 1728 349 1770 359
rect 1728 315 1736 349
rect 1728 299 1770 315
rect 1804 485 1870 493
rect 1804 451 1820 485
rect 1854 451 1870 485
rect 2143 485 2185 527
rect 2143 466 2151 485
rect 1804 417 1870 451
rect 1804 383 1820 417
rect 1854 383 1870 417
rect 1804 349 1870 383
rect 2011 451 2151 466
rect 2011 448 2185 451
rect 2011 385 2024 448
rect 2078 417 2185 448
rect 2078 385 2151 417
rect 2011 383 2151 385
rect 2011 359 2185 383
rect 1804 315 1820 349
rect 1854 315 1870 349
rect 1804 297 1870 315
rect 2143 349 2185 359
rect 2143 315 2151 349
rect 2143 299 2185 315
rect 2219 485 2285 493
rect 2219 451 2235 485
rect 2269 451 2285 485
rect 2558 485 2600 527
rect 2558 466 2566 485
rect 2219 417 2285 451
rect 2219 383 2235 417
rect 2269 383 2285 417
rect 2219 349 2285 383
rect 2426 451 2566 466
rect 2426 448 2600 451
rect 2426 385 2439 448
rect 2493 417 2600 448
rect 2493 385 2566 417
rect 2426 383 2566 385
rect 2426 359 2600 383
rect 2219 315 2235 349
rect 2269 315 2285 349
rect 2219 297 2285 315
rect 2558 349 2600 359
rect 2558 315 2566 349
rect 2558 299 2600 315
rect 2634 485 2700 493
rect 2634 451 2650 485
rect 2684 451 2700 485
rect 2634 417 2700 451
rect 2634 383 2650 417
rect 2684 383 2700 417
rect 2634 349 2700 383
rect 2634 315 2650 349
rect 2684 315 2700 349
rect 2634 297 2700 315
rect 164 263 210 297
rect 579 263 625 297
rect 994 263 1040 297
rect 1409 263 1455 297
rect 1824 263 1870 297
rect 2239 263 2285 297
rect 2654 263 2700 297
rect 2747 263 2795 289
rect -238 249 130 263
rect -238 215 80 249
rect 114 215 130 249
rect 164 249 545 263
rect 164 215 495 249
rect 529 215 545 249
rect 579 249 960 263
rect 579 215 910 249
rect 944 215 960 249
rect 994 249 1375 263
rect 994 215 1325 249
rect 1359 215 1375 249
rect 1409 249 1790 263
rect 1409 215 1740 249
rect 1774 215 1790 249
rect 1824 249 2205 263
rect 1824 215 2155 249
rect 2189 215 2205 249
rect 2239 249 2620 263
rect 2239 215 2570 249
rect 2604 215 2620 249
rect 2654 215 2926 263
rect -234 -128 -186 215
rect -64 165 110 181
rect 164 177 210 215
rect -64 160 76 165
rect -64 81 -51 160
rect 1 131 76 160
rect 1 97 110 131
rect 1 81 76 97
rect -64 63 76 81
rect -64 62 110 63
rect 64 17 110 62
rect 144 165 210 177
rect 144 131 160 165
rect 194 131 210 165
rect 144 97 210 131
rect 144 63 160 97
rect 194 63 210 97
rect 144 51 210 63
rect 351 165 525 181
rect 579 177 625 215
rect 351 160 491 165
rect 351 81 364 160
rect 416 131 491 160
rect 416 97 525 131
rect 416 81 491 97
rect 351 63 491 81
rect 351 62 525 63
rect 479 17 525 62
rect 559 165 625 177
rect 559 131 575 165
rect 609 131 625 165
rect 559 97 625 131
rect 559 63 575 97
rect 609 63 625 97
rect 559 51 625 63
rect 766 165 940 181
rect 994 177 1040 215
rect 766 160 906 165
rect 766 81 779 160
rect 831 131 906 160
rect 831 97 940 131
rect 831 81 906 97
rect 766 63 906 81
rect 766 62 940 63
rect 894 17 940 62
rect 974 165 1040 177
rect 974 131 990 165
rect 1024 131 1040 165
rect 974 97 1040 131
rect 974 63 990 97
rect 1024 63 1040 97
rect 974 51 1040 63
rect 1181 165 1355 181
rect 1409 177 1455 215
rect 1181 160 1321 165
rect 1181 81 1194 160
rect 1246 131 1321 160
rect 1246 97 1355 131
rect 1246 81 1321 97
rect 1181 63 1321 81
rect 1181 62 1355 63
rect 1309 17 1355 62
rect 1389 165 1455 177
rect 1389 131 1405 165
rect 1439 131 1455 165
rect 1389 97 1455 131
rect 1389 63 1405 97
rect 1439 63 1455 97
rect 1389 51 1455 63
rect 1596 165 1770 181
rect 1824 177 1870 215
rect 1596 160 1736 165
rect 1596 81 1609 160
rect 1661 131 1736 160
rect 1661 97 1770 131
rect 1661 81 1736 97
rect 1596 63 1736 81
rect 1596 62 1770 63
rect 1724 17 1770 62
rect 1804 165 1870 177
rect 1804 131 1820 165
rect 1854 131 1870 165
rect 1804 97 1870 131
rect 1804 63 1820 97
rect 1854 63 1870 97
rect 1804 51 1870 63
rect 2011 165 2185 181
rect 2239 177 2285 215
rect 2011 160 2151 165
rect 2011 81 2024 160
rect 2076 131 2151 160
rect 2076 97 2185 131
rect 2076 81 2151 97
rect 2011 63 2151 81
rect 2011 62 2185 63
rect 2139 17 2185 62
rect 2219 165 2285 177
rect 2219 131 2235 165
rect 2269 131 2285 165
rect 2219 97 2285 131
rect 2219 63 2235 97
rect 2269 63 2285 97
rect 2219 51 2285 63
rect 2426 165 2600 181
rect 2654 177 2700 215
rect 2426 160 2566 165
rect 2426 81 2439 160
rect 2491 131 2566 160
rect 2491 97 2600 131
rect 2491 81 2566 97
rect 2426 63 2566 81
rect 2426 62 2600 63
rect 2554 17 2600 62
rect 2634 165 2700 177
rect 2634 131 2650 165
rect 2684 131 2700 165
rect 2634 97 2700 131
rect 2634 63 2650 97
rect 2684 63 2700 97
rect 2634 51 2700 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
rect 415 -17 444 17
rect 478 -17 536 17
rect 570 -17 628 17
rect 662 -17 691 17
rect 830 -17 859 17
rect 893 -17 951 17
rect 985 -17 1043 17
rect 1077 -17 1106 17
rect 1245 -17 1274 17
rect 1308 -17 1366 17
rect 1400 -17 1458 17
rect 1492 -17 1521 17
rect 1660 -17 1689 17
rect 1723 -17 1781 17
rect 1815 -17 1873 17
rect 1907 -17 1936 17
rect 2075 -17 2104 17
rect 2138 -17 2196 17
rect 2230 -17 2288 17
rect 2322 -17 2351 17
rect 2490 -17 2519 17
rect 2553 -17 2611 17
rect 2645 -17 2703 17
rect 2737 -17 2766 17
rect 2878 -128 2926 215
rect -234 -176 2926 -128
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 444 527 478 561
rect 536 527 570 561
rect 628 527 662 561
rect 859 527 893 561
rect 951 527 985 561
rect 1043 527 1077 561
rect 1274 527 1308 561
rect 1366 527 1400 561
rect 1458 527 1492 561
rect 1689 527 1723 561
rect 1781 527 1815 561
rect 1873 527 1907 561
rect 2104 527 2138 561
rect 2196 527 2230 561
rect 2288 527 2322 561
rect 2519 527 2553 561
rect 2611 527 2645 561
rect 2703 527 2737 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 444 -17 478 17
rect 536 -17 570 17
rect 628 -17 662 17
rect 859 -17 893 17
rect 951 -17 985 17
rect 1043 -17 1077 17
rect 1274 -17 1308 17
rect 1366 -17 1400 17
rect 1458 -17 1492 17
rect 1689 -17 1723 17
rect 1781 -17 1815 17
rect 1873 -17 1907 17
rect 2104 -17 2138 17
rect 2196 -17 2230 17
rect 2288 -17 2322 17
rect 2519 -17 2553 17
rect 2611 -17 2645 17
rect 2703 -17 2737 17
<< metal1 >>
rect -69 592 -21 593
rect -101 561 2804 592
rect -101 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 444 561
rect 478 527 536 561
rect 570 527 628 561
rect 662 527 859 561
rect 893 527 951 561
rect 985 527 1043 561
rect 1077 527 1274 561
rect 1308 527 1366 561
rect 1400 527 1458 561
rect 1492 527 1689 561
rect 1723 527 1781 561
rect 1815 527 1873 561
rect 1907 527 2104 561
rect 2138 527 2196 561
rect 2230 527 2288 561
rect 2322 527 2519 561
rect 2553 527 2611 561
rect 2645 527 2703 561
rect 2737 527 2804 561
rect -101 496 2804 527
rect -101 17 2804 48
rect -101 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 444 17
rect 478 -17 536 17
rect 570 -17 628 17
rect 662 -17 859 17
rect 893 -17 951 17
rect 985 -17 1043 17
rect 1077 -17 1274 17
rect 1308 -17 1366 17
rect 1400 -17 1458 17
rect 1492 -17 1689 17
rect 1723 -17 1781 17
rect 1815 -17 1873 17
rect 1907 -17 2104 17
rect 2138 -17 2196 17
rect 2230 -17 2288 17
rect 2322 -17 2519 17
rect 2553 -17 2611 17
rect 2645 -17 2703 17
rect 2737 -17 2804 17
rect -101 -48 2804 -17
<< labels >>
flabel metal1 -69 545 -21 593 1 FreeSans 400 0 0 0 VDD
port 2 n
flabel metal1 -65 -10 -17 38 1 FreeSans 400 0 0 0 gnd
port 3 n
flabel locali 2747 241 2795 289 1 FreeSans 400 0 0 0 out
port 1 n
flabel locali 72 221 106 255 0 FreeSans 340 0 0 0 inv1_0[0].A
flabel locali 164 289 198 323 0 FreeSans 340 0 0 0 inv1_0[0].Y
flabel metal1 29 527 63 561 0 FreeSans 200 0 0 0 inv1_0[0].VPWR
flabel metal1 29 -17 63 17 0 FreeSans 200 0 0 0 inv1_0[0].VGND
rlabel comment 0 0 0 0 4 inv1_0[0].inv_1
flabel locali 487 221 521 255 0 FreeSans 340 0 0 0 inv1_0[1].A
flabel locali 579 289 613 323 0 FreeSans 340 0 0 0 inv1_0[1].Y
flabel metal1 444 527 478 561 0 FreeSans 200 0 0 0 inv1_0[1].VPWR
flabel metal1 444 -17 478 17 0 FreeSans 200 0 0 0 inv1_0[1].VGND
rlabel comment 415 0 415 0 4 inv1_0[1].inv_1
flabel locali 902 221 936 255 0 FreeSans 340 0 0 0 inv1_0[2].A
flabel locali 994 289 1028 323 0 FreeSans 340 0 0 0 inv1_0[2].Y
flabel metal1 859 527 893 561 0 FreeSans 200 0 0 0 inv1_0[2].VPWR
flabel metal1 859 -17 893 17 0 FreeSans 200 0 0 0 inv1_0[2].VGND
rlabel comment 830 0 830 0 4 inv1_0[2].inv_1
flabel locali 1317 221 1351 255 0 FreeSans 340 0 0 0 inv1_0[3].A
flabel locali 1409 289 1443 323 0 FreeSans 340 0 0 0 inv1_0[3].Y
flabel metal1 1274 527 1308 561 0 FreeSans 200 0 0 0 inv1_0[3].VPWR
flabel metal1 1274 -17 1308 17 0 FreeSans 200 0 0 0 inv1_0[3].VGND
rlabel comment 1245 0 1245 0 4 inv1_0[3].inv_1
flabel locali 1732 221 1766 255 0 FreeSans 340 0 0 0 inv1_0[4].A
flabel locali 1824 289 1858 323 0 FreeSans 340 0 0 0 inv1_0[4].Y
flabel metal1 1689 527 1723 561 0 FreeSans 200 0 0 0 inv1_0[4].VPWR
flabel metal1 1689 -17 1723 17 0 FreeSans 200 0 0 0 inv1_0[4].VGND
rlabel comment 1660 0 1660 0 4 inv1_0[4].inv_1
flabel locali 2147 221 2181 255 0 FreeSans 340 0 0 0 inv1_0[5].A
flabel locali 2239 289 2273 323 0 FreeSans 340 0 0 0 inv1_0[5].Y
flabel metal1 2104 527 2138 561 0 FreeSans 200 0 0 0 inv1_0[5].VPWR
flabel metal1 2104 -17 2138 17 0 FreeSans 200 0 0 0 inv1_0[5].VGND
rlabel comment 2075 0 2075 0 4 inv1_0[5].inv_1
flabel locali 2562 221 2596 255 0 FreeSans 340 0 0 0 inv1_0[6].A
flabel locali 2654 289 2688 323 0 FreeSans 340 0 0 0 inv1_0[6].Y
flabel metal1 2519 527 2553 561 0 FreeSans 200 0 0 0 inv1_0[6].VPWR
flabel metal1 2519 -17 2553 17 0 FreeSans 200 0 0 0 inv1_0[6].VGND
rlabel comment 2490 0 2490 0 4 inv1_0[6].inv_1
<< end >>
