magic
tech sky130A
magscale 1 2
timestamp 1608329073
<< locali >>
rect -214 217 -65 265
rect 1090 217 1264 265
rect -214 -56 -166 217
rect 1216 -56 1264 217
rect -214 -104 1264 -56
<< metal1 >>
rect -95 508 -23 577
rect -91 -32 -28 33
use inv1  inv1_0 layout
array 0 2 415 0 0 640
timestamp 1608267076
transform 1 0 -6 0 1 2
box -101 -48 314 592
<< labels >>
flabel locali 1173 225 1233 256 1 FreeSans 400 0 0 0 out
port 1 n
flabel metal1 -95 508 -23 577 1 FreeSans 400 0 0 0 vdd
port 3 n
flabel metal1 -91 -32 -28 33 1 FreeSans 400 0 0 0 gnd
port 2 n
<< end >>
