* Simple inverter

.subckt inv1 A VGND VNB VPB VPWR Y

X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u

.ends
