* Simple inverter

.subckt inv1 A Y VPWR VGND

X0 Y A VGND VGND sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 Y A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u

.ends
* Ring oscillator circuit

.subckt ringosc out vdd gnd

X0 out y1 vdd gnd inv1
X1 y1 y2 vdd gnd inv1
X2 y2 y3 vdd gnd inv1
X3 y3 y4 vdd gnd inv1
X4 y4 y5 vdd gnd inv1
X5 y5 y6 vdd gnd inv1
X6 y6 out vdd gnd inv1


.ends
