magic
tech sky130A
magscale 1 2
timestamp 1608267076
<< nwell >>
rect -101 261 314 582
<< pwell >>
rect 29 -17 63 17
<< scnmos >>
rect 120 47 150 177
<< scpmoshvt >>
rect 120 297 150 497
<< ndiff >>
rect 68 165 120 177
rect 68 131 76 165
rect 110 131 120 165
rect 68 97 120 131
rect 68 63 76 97
rect 110 63 120 97
rect 68 47 120 63
rect 150 165 202 177
rect 150 131 160 165
rect 194 131 202 165
rect 150 97 202 131
rect 150 63 160 97
rect 194 63 202 97
rect 150 47 202 63
<< pdiff >>
rect 68 485 120 497
rect 68 451 76 485
rect 110 451 120 485
rect 68 417 120 451
rect 68 383 76 417
rect 110 383 120 417
rect 68 349 120 383
rect 68 315 76 349
rect 110 315 120 349
rect 68 297 120 315
rect 150 485 202 497
rect 150 451 160 485
rect 194 451 202 485
rect 150 417 202 451
rect 150 383 160 417
rect 194 383 202 417
rect 150 349 202 383
rect 150 315 160 349
rect 194 315 202 349
rect 150 297 202 315
<< ndiffc >>
rect 76 131 110 165
rect 76 63 110 97
rect 160 131 194 165
rect 160 63 194 97
<< pdiffc >>
rect 76 451 110 485
rect 76 383 110 417
rect 76 315 110 349
rect 160 451 194 485
rect 160 383 194 417
rect 160 315 194 349
<< psubdiff >>
rect -64 160 14 190
rect -64 81 -51 160
rect 1 81 14 160
rect -64 55 14 81
<< nsubdiff >>
rect -64 448 14 479
rect -64 385 -51 448
rect 3 385 14 448
rect -64 336 14 385
<< psubdiffcont >>
rect -51 81 1 160
<< nsubdiffcont >>
rect -51 385 3 448
<< poly >>
rect 120 497 150 523
rect 120 265 150 297
rect 64 249 150 265
rect 64 215 80 249
rect 114 215 150 249
rect 64 199 150 215
rect 120 177 150 199
rect 120 21 150 47
<< polycont >>
rect 80 215 114 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 68 485 110 527
rect 68 466 76 485
rect -64 451 76 466
rect -64 448 110 451
rect -64 385 -51 448
rect 3 417 110 448
rect 3 385 76 417
rect -64 383 76 385
rect -64 359 110 383
rect 68 349 110 359
rect 68 315 76 349
rect 68 299 110 315
rect 144 485 210 493
rect 144 451 160 485
rect 194 451 210 485
rect 144 417 210 451
rect 144 383 160 417
rect 194 383 210 417
rect 144 349 210 383
rect 144 315 160 349
rect 194 315 210 349
rect 144 297 210 315
rect 164 263 210 297
rect -101 249 130 263
rect -101 215 80 249
rect 114 215 130 249
rect 164 215 314 263
rect -64 165 110 181
rect 164 177 210 215
rect -64 160 76 165
rect -64 81 -51 160
rect 1 131 76 160
rect 1 97 110 131
rect 1 81 76 97
rect -64 63 76 81
rect -64 62 110 63
rect 64 17 110 62
rect 144 165 210 177
rect 144 131 160 165
rect 194 131 210 165
rect 144 97 210 131
rect 144 63 160 97
rect 194 63 210 97
rect 144 51 210 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
<< metal1 >>
rect -101 561 314 592
rect -101 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 314 561
rect -101 496 314 527
rect -101 17 314 48
rect -101 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 314 17
rect -101 -48 314 -17
<< labels >>
flabel locali s 164 289 198 323 0 FreeSans 340 0 0 0 Y
port 1 nsew
flabel locali s 72 221 106 255 0 FreeSans 340 0 0 0 A
port 2 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 4 nsew
rlabel comment s 0 0 0 0 4 inv_1
<< properties >>
string FIXED_BBOX 0 0 276 544
string path 0.000 0.000 1.380 0.000 
<< end >>
