* Include SKY130 libraries
.lib "/path/to/skywater-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice" tt
