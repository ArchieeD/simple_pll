* Testbench for a ring oscillator

* YOUR IMPLEMENTATION HERE
X0 ro_out vddi 0 ringosc
X1 ro_out 0 0 vddo vddo out

V0 vddi 0 0.65
V1 vddo 0 0.80

.nodeset V(ro_out)=0
